/*-----------------------------------------------------------------------------*/
/*  Common header for saxi2maxi.v                                              */
/*-----------------------------------------------------------------------------*/

//`define			BUFG_ENABLE
`define			CPU_RESET_CNT			32'h0010_0000		// Min=32'h0000_0010,Max=32'hFFFF_FFFE
`define			USER_RESET_CNT			32'h0100_0000		// Min=32'h0000_0010,Max=32'hFFFF_FFFE
`define			PERI_RESET_CNT			32'h0200_0000		// Min=32'h0000_0010,Max=32'hFFFF_FFFE



